//ram
//バス幅2048bit
module ram (
    input clk_h,    // Clock
    input clk_l,    // Clock(負論理)
    input w_e, // Write Enable
    //input rst_n,  // Asynchronous reset active low
    input  wire [15:0]read_adr,   //アドレスバス
    input  wire [15:0]write_adr,   //アドレスバス
    output reg  [1023:0]read_data, //メモリからのデータ出力
    input  wire [1023:0]write_data //メモリへ書き込むデータ入力
);

reg [131072:0]ram;

always @(posedge clk_h or negedge clk_l) begin
    read_data <= {ram[read_adr+1023],ram[read_adr+1022],ram[read_adr+1021],ram[read_adr+1020],ram[read_adr+1019],ram[read_adr+1018],ram[read_adr+1017],ram[read_adr+1016],ram[read_adr+1015],ram[read_adr+1014],ram[read_adr+1013],ram[read_adr+1012],ram[read_adr+1011],ram[read_adr+1010],ram[read_adr+1009],ram[read_adr+1008],ram[read_adr+1007],ram[read_adr+1006],ram[read_adr+1005],ram[read_adr+1004],ram[read_adr+1003],ram[read_adr+1002],ram[read_adr+1001],ram[read_adr+1000],ram[read_adr+999],ram[read_adr+998],ram[read_adr+997],ram[read_adr+996],ram[read_adr+995],ram[read_adr+994],ram[read_adr+993],ram[read_adr+992],ram[read_adr+991],ram[read_adr+990],ram[read_adr+989],ram[read_adr+988],ram[read_adr+987],ram[read_adr+986],ram[read_adr+985],ram[read_adr+984],ram[read_adr+983],ram[read_adr+982],ram[read_adr+981],ram[read_adr+980],ram[read_adr+979],ram[read_adr+978],ram[read_adr+977],ram[read_adr+976],ram[read_adr+975],ram[read_adr+974],ram[read_adr+973],ram[read_adr+972],ram[read_adr+971],ram[read_adr+970],ram[read_adr+969],ram[read_adr+968],ram[read_adr+967],ram[read_adr+966],ram[read_adr+965],ram[read_adr+964],ram[read_adr+963],ram[read_adr+962],ram[read_adr+961],ram[read_adr+960],ram[read_adr+959],ram[read_adr+958],ram[read_adr+957],ram[read_adr+956],ram[read_adr+955],ram[read_adr+954],ram[read_adr+953],ram[read_adr+952],ram[read_adr+951],ram[read_adr+950],ram[read_adr+949],ram[read_adr+948],ram[read_adr+947],ram[read_adr+946],ram[read_adr+945],ram[read_adr+944],ram[read_adr+943],ram[read_adr+942],ram[read_adr+941],ram[read_adr+940],ram[read_adr+939],ram[read_adr+938],ram[read_adr+937],ram[read_adr+936],ram[read_adr+935],ram[read_adr+934],ram[read_adr+933],ram[read_adr+932],ram[read_adr+931],ram[read_adr+930],ram[read_adr+929],ram[read_adr+928],ram[read_adr+927],ram[read_adr+926],ram[read_adr+925],ram[read_adr+924],ram[read_adr+923],ram[read_adr+922],ram[read_adr+921],ram[read_adr+920],ram[read_adr+919],ram[read_adr+918],ram[read_adr+917],ram[read_adr+916],ram[read_adr+915],ram[read_adr+914],ram[read_adr+913],ram[read_adr+912],ram[read_adr+911],ram[read_adr+910],ram[read_adr+909],ram[read_adr+908],ram[read_adr+907],ram[read_adr+906],ram[read_adr+905],ram[read_adr+904],ram[read_adr+903],ram[read_adr+902],ram[read_adr+901],ram[read_adr+900],ram[read_adr+899],ram[read_adr+898],ram[read_adr+897],ram[read_adr+896],ram[read_adr+895],ram[read_adr+894],ram[read_adr+893],ram[read_adr+892],ram[read_adr+891],ram[read_adr+890],ram[read_adr+889],ram[read_adr+888],ram[read_adr+887],ram[read_adr+886],ram[read_adr+885],ram[read_adr+884],ram[read_adr+883],ram[read_adr+882],ram[read_adr+881],ram[read_adr+880],ram[read_adr+879],ram[read_adr+878],ram[read_adr+877],ram[read_adr+876],ram[read_adr+875],ram[read_adr+874],ram[read_adr+873],ram[read_adr+872],ram[read_adr+871],ram[read_adr+870],ram[read_adr+869],ram[read_adr+868],ram[read_adr+867],ram[read_adr+866],ram[read_adr+865],ram[read_adr+864],ram[read_adr+863],ram[read_adr+862],ram[read_adr+861],ram[read_adr+860],ram[read_adr+859],ram[read_adr+858],ram[read_adr+857],ram[read_adr+856],ram[read_adr+855],ram[read_adr+854],ram[read_adr+853],ram[read_adr+852],ram[read_adr+851],ram[read_adr+850],ram[read_adr+849],ram[read_adr+848],ram[read_adr+847],ram[read_adr+846],ram[read_adr+845],ram[read_adr+844],ram[read_adr+843],ram[read_adr+842],ram[read_adr+841],ram[read_adr+840],ram[read_adr+839],ram[read_adr+838],ram[read_adr+837],ram[read_adr+836],ram[read_adr+835],ram[read_adr+834],ram[read_adr+833],ram[read_adr+832],ram[read_adr+831],ram[read_adr+830],ram[read_adr+829],ram[read_adr+828],ram[read_adr+827],ram[read_adr+826],ram[read_adr+825],ram[read_adr+824],ram[read_adr+823],ram[read_adr+822],ram[read_adr+821],ram[read_adr+820],ram[read_adr+819],ram[read_adr+818],ram[read_adr+817],ram[read_adr+816],ram[read_adr+815],ram[read_adr+814],ram[read_adr+813],ram[read_adr+812],ram[read_adr+811],ram[read_adr+810],ram[read_adr+809],ram[read_adr+808],ram[read_adr+807],ram[read_adr+806],ram[read_adr+805],ram[read_adr+804],ram[read_adr+803],ram[read_adr+802],ram[read_adr+801],ram[read_adr+800],ram[read_adr+799],ram[read_adr+798],ram[read_adr+797],ram[read_adr+796],ram[read_adr+795],ram[read_adr+794],ram[read_adr+793],ram[read_adr+792],ram[read_adr+791],ram[read_adr+790],ram[read_adr+789],ram[read_adr+788],ram[read_adr+787],ram[read_adr+786],ram[read_adr+785],ram[read_adr+784],ram[read_adr+783],ram[read_adr+782],ram[read_adr+781],ram[read_adr+780],ram[read_adr+779],ram[read_adr+778],ram[read_adr+777],ram[read_adr+776],ram[read_adr+775],ram[read_adr+774],ram[read_adr+773],ram[read_adr+772],ram[read_adr+771],ram[read_adr+770],ram[read_adr+769],ram[read_adr+768],ram[read_adr+767],ram[read_adr+766],ram[read_adr+765],ram[read_adr+764],ram[read_adr+763],ram[read_adr+762],ram[read_adr+761],ram[read_adr+760],ram[read_adr+759],ram[read_adr+758],ram[read_adr+757],ram[read_adr+756],ram[read_adr+755],ram[read_adr+754],ram[read_adr+753],ram[read_adr+752],ram[read_adr+751],ram[read_adr+750],ram[read_adr+749],ram[read_adr+748],ram[read_adr+747],ram[read_adr+746],ram[read_adr+745],ram[read_adr+744],ram[read_adr+743],ram[read_adr+742],ram[read_adr+741],ram[read_adr+740],ram[read_adr+739],ram[read_adr+738],ram[read_adr+737],ram[read_adr+736],ram[read_adr+735],ram[read_adr+734],ram[read_adr+733],ram[read_adr+732],ram[read_adr+731],ram[read_adr+730],ram[read_adr+729],ram[read_adr+728],ram[read_adr+727],ram[read_adr+726],ram[read_adr+725],ram[read_adr+724],ram[read_adr+723],ram[read_adr+722],ram[read_adr+721],ram[read_adr+720],ram[read_adr+719],ram[read_adr+718],ram[read_adr+717],ram[read_adr+716],ram[read_adr+715],ram[read_adr+714],ram[read_adr+713],ram[read_adr+712],ram[read_adr+711],ram[read_adr+710],ram[read_adr+709],ram[read_adr+708],ram[read_adr+707],ram[read_adr+706],ram[read_adr+705],ram[read_adr+704],ram[read_adr+703],ram[read_adr+702],ram[read_adr+701],ram[read_adr+700],ram[read_adr+699],ram[read_adr+698],ram[read_adr+697],ram[read_adr+696],ram[read_adr+695],ram[read_adr+694],ram[read_adr+693],ram[read_adr+692],ram[read_adr+691],ram[read_adr+690],ram[read_adr+689],ram[read_adr+688],ram[read_adr+687],ram[read_adr+686],ram[read_adr+685],ram[read_adr+684],ram[read_adr+683],ram[read_adr+682],ram[read_adr+681],ram[read_adr+680],ram[read_adr+679],ram[read_adr+678],ram[read_adr+677],ram[read_adr+676],ram[read_adr+675],ram[read_adr+674],ram[read_adr+673],ram[read_adr+672],ram[read_adr+671],ram[read_adr+670],ram[read_adr+669],ram[read_adr+668],ram[read_adr+667],ram[read_adr+666],ram[read_adr+665],ram[read_adr+664],ram[read_adr+663],ram[read_adr+662],ram[read_adr+661],ram[read_adr+660],ram[read_adr+659],ram[read_adr+658],ram[read_adr+657],ram[read_adr+656],ram[read_adr+655],ram[read_adr+654],ram[read_adr+653],ram[read_adr+652],ram[read_adr+651],ram[read_adr+650],ram[read_adr+649],ram[read_adr+648],ram[read_adr+647],ram[read_adr+646],ram[read_adr+645],ram[read_adr+644],ram[read_adr+643],ram[read_adr+642],ram[read_adr+641],ram[read_adr+640],ram[read_adr+639],ram[read_adr+638],ram[read_adr+637],ram[read_adr+636],ram[read_adr+635],ram[read_adr+634],ram[read_adr+633],ram[read_adr+632],ram[read_adr+631],ram[read_adr+630],ram[read_adr+629],ram[read_adr+628],ram[read_adr+627],ram[read_adr+626],ram[read_adr+625],ram[read_adr+624],ram[read_adr+623],ram[read_adr+622],ram[read_adr+621],ram[read_adr+620],ram[read_adr+619],ram[read_adr+618],ram[read_adr+617],ram[read_adr+616],ram[read_adr+615],ram[read_adr+614],ram[read_adr+613],ram[read_adr+612],ram[read_adr+611],ram[read_adr+610],ram[read_adr+609],ram[read_adr+608],ram[read_adr+607],ram[read_adr+606],ram[read_adr+605],ram[read_adr+604],ram[read_adr+603],ram[read_adr+602],ram[read_adr+601],ram[read_adr+600],ram[read_adr+599],ram[read_adr+598],ram[read_adr+597],ram[read_adr+596],ram[read_adr+595],ram[read_adr+594],ram[read_adr+593],ram[read_adr+592],ram[read_adr+591],ram[read_adr+590],ram[read_adr+589],ram[read_adr+588],ram[read_adr+587],ram[read_adr+586],ram[read_adr+585],ram[read_adr+584],ram[read_adr+583],ram[read_adr+582],ram[read_adr+581],ram[read_adr+580],ram[read_adr+579],ram[read_adr+578],ram[read_adr+577],ram[read_adr+576],ram[read_adr+575],ram[read_adr+574],ram[read_adr+573],ram[read_adr+572],ram[read_adr+571],ram[read_adr+570],ram[read_adr+569],ram[read_adr+568],ram[read_adr+567],ram[read_adr+566],ram[read_adr+565],ram[read_adr+564],ram[read_adr+563],ram[read_adr+562],ram[read_adr+561],ram[read_adr+560],ram[read_adr+559],ram[read_adr+558],ram[read_adr+557],ram[read_adr+556],ram[read_adr+555],ram[read_adr+554],ram[read_adr+553],ram[read_adr+552],ram[read_adr+551],ram[read_adr+550],ram[read_adr+549],ram[read_adr+548],ram[read_adr+547],ram[read_adr+546],ram[read_adr+545],ram[read_adr+544],ram[read_adr+543],ram[read_adr+542],ram[read_adr+541],ram[read_adr+540],ram[read_adr+539],ram[read_adr+538],ram[read_adr+537],ram[read_adr+536],ram[read_adr+535],ram[read_adr+534],ram[read_adr+533],ram[read_adr+532],ram[read_adr+531],ram[read_adr+530],ram[read_adr+529],ram[read_adr+528],ram[read_adr+527],ram[read_adr+526],ram[read_adr+525],ram[read_adr+524],ram[read_adr+523],ram[read_adr+522],ram[read_adr+521],ram[read_adr+520],ram[read_adr+519],ram[read_adr+518],ram[read_adr+517],ram[read_adr+516],ram[read_adr+515],ram[read_adr+514],ram[read_adr+513],ram[read_adr+512],ram[read_adr+511],ram[read_adr+510],ram[read_adr+509],ram[read_adr+508],ram[read_adr+507],ram[read_adr+506],ram[read_adr+505],ram[read_adr+504],ram[read_adr+503],ram[read_adr+502],ram[read_adr+501],ram[read_adr+500],ram[read_adr+499],ram[read_adr+498],ram[read_adr+497],ram[read_adr+496],ram[read_adr+495],ram[read_adr+494],ram[read_adr+493],ram[read_adr+492],ram[read_adr+491],ram[read_adr+490],ram[read_adr+489],ram[read_adr+488],ram[read_adr+487],ram[read_adr+486],ram[read_adr+485],ram[read_adr+484],ram[read_adr+483],ram[read_adr+482],ram[read_adr+481],ram[read_adr+480],ram[read_adr+479],ram[read_adr+478],ram[read_adr+477],ram[read_adr+476],ram[read_adr+475],ram[read_adr+474],ram[read_adr+473],ram[read_adr+472],ram[read_adr+471],ram[read_adr+470],ram[read_adr+469],ram[read_adr+468],ram[read_adr+467],ram[read_adr+466],ram[read_adr+465],ram[read_adr+464],ram[read_adr+463],ram[read_adr+462],ram[read_adr+461],ram[read_adr+460],ram[read_adr+459],ram[read_adr+458],ram[read_adr+457],ram[read_adr+456],ram[read_adr+455],ram[read_adr+454],ram[read_adr+453],ram[read_adr+452],ram[read_adr+451],ram[read_adr+450],ram[read_adr+449],ram[read_adr+448],ram[read_adr+447],ram[read_adr+446],ram[read_adr+445],ram[read_adr+444],ram[read_adr+443],ram[read_adr+442],ram[read_adr+441],ram[read_adr+440],ram[read_adr+439],ram[read_adr+438],ram[read_adr+437],ram[read_adr+436],ram[read_adr+435],ram[read_adr+434],ram[read_adr+433],ram[read_adr+432],ram[read_adr+431],ram[read_adr+430],ram[read_adr+429],ram[read_adr+428],ram[read_adr+427],ram[read_adr+426],ram[read_adr+425],ram[read_adr+424],ram[read_adr+423],ram[read_adr+422],ram[read_adr+421],ram[read_adr+420],ram[read_adr+419],ram[read_adr+418],ram[read_adr+417],ram[read_adr+416],ram[read_adr+415],ram[read_adr+414],ram[read_adr+413],ram[read_adr+412],ram[read_adr+411],ram[read_adr+410],ram[read_adr+409],ram[read_adr+408],ram[read_adr+407],ram[read_adr+406],ram[read_adr+405],ram[read_adr+404],ram[read_adr+403],ram[read_adr+402],ram[read_adr+401],ram[read_adr+400],ram[read_adr+399],ram[read_adr+398],ram[read_adr+397],ram[read_adr+396],ram[read_adr+395],ram[read_adr+394],ram[read_adr+393],ram[read_adr+392],ram[read_adr+391],ram[read_adr+390],ram[read_adr+389],ram[read_adr+388],ram[read_adr+387],ram[read_adr+386],ram[read_adr+385],ram[read_adr+384],ram[read_adr+383],ram[read_adr+382],ram[read_adr+381],ram[read_adr+380],ram[read_adr+379],ram[read_adr+378],ram[read_adr+377],ram[read_adr+376],ram[read_adr+375],ram[read_adr+374],ram[read_adr+373],ram[read_adr+372],ram[read_adr+371],ram[read_adr+370],ram[read_adr+369],ram[read_adr+368],ram[read_adr+367],ram[read_adr+366],ram[read_adr+365],ram[read_adr+364],ram[read_adr+363],ram[read_adr+362],ram[read_adr+361],ram[read_adr+360],ram[read_adr+359],ram[read_adr+358],ram[read_adr+357],ram[read_adr+356],ram[read_adr+355],ram[read_adr+354],ram[read_adr+353],ram[read_adr+352],ram[read_adr+351],ram[read_adr+350],ram[read_adr+349],ram[read_adr+348],ram[read_adr+347],ram[read_adr+346],ram[read_adr+345],ram[read_adr+344],ram[read_adr+343],ram[read_adr+342],ram[read_adr+341],ram[read_adr+340],ram[read_adr+339],ram[read_adr+338],ram[read_adr+337],ram[read_adr+336],ram[read_adr+335],ram[read_adr+334],ram[read_adr+333],ram[read_adr+332],ram[read_adr+331],ram[read_adr+330],ram[read_adr+329],ram[read_adr+328],ram[read_adr+327],ram[read_adr+326],ram[read_adr+325],ram[read_adr+324],ram[read_adr+323],ram[read_adr+322],ram[read_adr+321],ram[read_adr+320],ram[read_adr+319],ram[read_adr+318],ram[read_adr+317],ram[read_adr+316],ram[read_adr+315],ram[read_adr+314],ram[read_adr+313],ram[read_adr+312],ram[read_adr+311],ram[read_adr+310],ram[read_adr+309],ram[read_adr+308],ram[read_adr+307],ram[read_adr+306],ram[read_adr+305],ram[read_adr+304],ram[read_adr+303],ram[read_adr+302],ram[read_adr+301],ram[read_adr+300],ram[read_adr+299],ram[read_adr+298],ram[read_adr+297],ram[read_adr+296],ram[read_adr+295],ram[read_adr+294],ram[read_adr+293],ram[read_adr+292],ram[read_adr+291],ram[read_adr+290],ram[read_adr+289],ram[read_adr+288],ram[read_adr+287],ram[read_adr+286],ram[read_adr+285],ram[read_adr+284],ram[read_adr+283],ram[read_adr+282],ram[read_adr+281],ram[read_adr+280],ram[read_adr+279],ram[read_adr+278],ram[read_adr+277],ram[read_adr+276],ram[read_adr+275],ram[read_adr+274],ram[read_adr+273],ram[read_adr+272],ram[read_adr+271],ram[read_adr+270],ram[read_adr+269],ram[read_adr+268],ram[read_adr+267],ram[read_adr+266],ram[read_adr+265],ram[read_adr+264],ram[read_adr+263],ram[read_adr+262],ram[read_adr+261],ram[read_adr+260],ram[read_adr+259],ram[read_adr+258],ram[read_adr+257],ram[read_adr+256],ram[read_adr+255],ram[read_adr+254],ram[read_adr+253],ram[read_adr+252],ram[read_adr+251],ram[read_adr+250],ram[read_adr+249],ram[read_adr+248],ram[read_adr+247],ram[read_adr+246],ram[read_adr+245],ram[read_adr+244],ram[read_adr+243],ram[read_adr+242],ram[read_adr+241],ram[read_adr+240],ram[read_adr+239],ram[read_adr+238],ram[read_adr+237],ram[read_adr+236],ram[read_adr+235],ram[read_adr+234],ram[read_adr+233],ram[read_adr+232],ram[read_adr+231],ram[read_adr+230],ram[read_adr+229],ram[read_adr+228],ram[read_adr+227],ram[read_adr+226],ram[read_adr+225],ram[read_adr+224],ram[read_adr+223],ram[read_adr+222],ram[read_adr+221],ram[read_adr+220],ram[read_adr+219],ram[read_adr+218],ram[read_adr+217],ram[read_adr+216],ram[read_adr+215],ram[read_adr+214],ram[read_adr+213],ram[read_adr+212],ram[read_adr+211],ram[read_adr+210],ram[read_adr+209],ram[read_adr+208],ram[read_adr+207],ram[read_adr+206],ram[read_adr+205],ram[read_adr+204],ram[read_adr+203],ram[read_adr+202],ram[read_adr+201],ram[read_adr+200],ram[read_adr+199],ram[read_adr+198],ram[read_adr+197],ram[read_adr+196],ram[read_adr+195],ram[read_adr+194],ram[read_adr+193],ram[read_adr+192],ram[read_adr+191],ram[read_adr+190],ram[read_adr+189],ram[read_adr+188],ram[read_adr+187],ram[read_adr+186],ram[read_adr+185],ram[read_adr+184],ram[read_adr+183],ram[read_adr+182],ram[read_adr+181],ram[read_adr+180],ram[read_adr+179],ram[read_adr+178],ram[read_adr+177],ram[read_adr+176],ram[read_adr+175],ram[read_adr+174],ram[read_adr+173],ram[read_adr+172],ram[read_adr+171],ram[read_adr+170],ram[read_adr+169],ram[read_adr+168],ram[read_adr+167],ram[read_adr+166],ram[read_adr+165],ram[read_adr+164],ram[read_adr+163],ram[read_adr+162],ram[read_adr+161],ram[read_adr+160],ram[read_adr+159],ram[read_adr+158],ram[read_adr+157],ram[read_adr+156],ram[read_adr+155],ram[read_adr+154],ram[read_adr+153],ram[read_adr+152],ram[read_adr+151],ram[read_adr+150],ram[read_adr+149],ram[read_adr+148],ram[read_adr+147],ram[read_adr+146],ram[read_adr+145],ram[read_adr+144],ram[read_adr+143],ram[read_adr+142],ram[read_adr+141],ram[read_adr+140],ram[read_adr+139],ram[read_adr+138],ram[read_adr+137],ram[read_adr+136],ram[read_adr+135],ram[read_adr+134],ram[read_adr+133],ram[read_adr+132],ram[read_adr+131],ram[read_adr+130],ram[read_adr+129],ram[read_adr+128],ram[read_adr+127],ram[read_adr+126],ram[read_adr+125],ram[read_adr+124],ram[read_adr+123],ram[read_adr+122],ram[read_adr+121],ram[read_adr+120],ram[read_adr+119],ram[read_adr+118],ram[read_adr+117],ram[read_adr+116],ram[read_adr+115],ram[read_adr+114],ram[read_adr+113],ram[read_adr+112],ram[read_adr+111],ram[read_adr+110],ram[read_adr+109],ram[read_adr+108],ram[read_adr+107],ram[read_adr+106],ram[read_adr+105],ram[read_adr+104],ram[read_adr+103],ram[read_adr+102],ram[read_adr+101],ram[read_adr+100],ram[read_adr+99],ram[read_adr+98],ram[read_adr+97],ram[read_adr+96],ram[read_adr+95],ram[read_adr+94],ram[read_adr+93],ram[read_adr+92],ram[read_adr+91],ram[read_adr+90],ram[read_adr+89],ram[read_adr+88],ram[read_adr+87],ram[read_adr+86],ram[read_adr+85],ram[read_adr+84],ram[read_adr+83],ram[read_adr+82],ram[read_adr+81],ram[read_adr+80],ram[read_adr+79],ram[read_adr+78],ram[read_adr+77],ram[read_adr+76],ram[read_adr+75],ram[read_adr+74],ram[read_adr+73],ram[read_adr+72],ram[read_adr+71],ram[read_adr+70],ram[read_adr+69],ram[read_adr+68],ram[read_adr+67],ram[read_adr+66],ram[read_adr+65],ram[read_adr+64],ram[read_adr+63],ram[read_adr+62],ram[read_adr+61],ram[read_adr+60],ram[read_adr+59],ram[read_adr+58],ram[read_adr+57],ram[read_adr+56],ram[read_adr+55],ram[read_adr+54],ram[read_adr+53],ram[read_adr+52],ram[read_adr+51],ram[read_adr+50],ram[read_adr+49],ram[read_adr+48],ram[read_adr+47],ram[read_adr+46],ram[read_adr+45],ram[read_adr+44],ram[read_adr+43],ram[read_adr+42],ram[read_adr+41],ram[read_adr+40],ram[read_adr+39],ram[read_adr+38],ram[read_adr+37],ram[read_adr+36],ram[read_adr+35],ram[read_adr+34],ram[read_adr+33],ram[read_adr+32],ram[read_adr+31],ram[read_adr+30],ram[read_adr+29],ram[read_adr+28],ram[read_adr+27],ram[read_adr+26],ram[read_adr+25],ram[read_adr+24],ram[read_adr+23],ram[read_adr+22],ram[read_adr+21],ram[read_adr+20],ram[read_adr+19],ram[read_adr+18],ram[read_adr+17],ram[read_adr+16],ram[read_adr+15],ram[read_adr+14],ram[read_adr+13],ram[read_adr+12],ram[read_adr+11],ram[read_adr+10],ram[read_adr+9],ram[read_adr+8],ram[read_adr+7],ram[read_adr+6],ram[read_adr+5],ram[read_adr+4],ram[read_adr+3],ram[read_adr+2],ram[read_adr+1],ram[read_adr+0]};
    //if(write_adr+i<4096)
        //ram[write_adr*8192:write_adr*8] <= write_data;
    //end
end

endmodule