module insdecoder (
    /*--------------------------------------------------*/
    input wire [1023:0]ins,//命令本体のinput
    /*--------------------------------------------------*/
    output wire meta_inst,//通常の演算命令かどうかの MSB
    output wire [6:0]eval_len, //評価する長さMSB-1~7bit
    output wire [15:0]operand,  //特殊命令へのオペランド(ジャンプ等) 残り16bit
    /*--------------------------------------------------*/
    output wire [7:0]alu_code, //ALUへのコード 8bit
    output wire [7:0]alu_src,  //ALUへのソース
    output wire [7:0]alu_dst,  //ALUへのデスティネーション
    /*--------------------------------------------------*/
    output wire [15:0]next
    /*--------------------------------------------------*/
);

/*--------------------------------------------------*/

/*--------------------------------------------------*/
endmodule